//Jtag+ tap con
